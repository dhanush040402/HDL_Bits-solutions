module top_module (
    input clk,
    input reset,
    input [31:0] in,
    output [31:0] out
);

    reg [31:0] i;	
  
  always @(posedge clk) begin
      i <= in;
      if(reset) 
        out <= 0;
      else begin
        out <= out | (i & ~in);
      end
  end
endmodule
